library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

package Imageqq is

	constant DIS_MAX_X :integer:= 80;		--横坐标
	constant DIS_MAX_Y :integer:= 60;		--纵坐标

	subtype MemVideoPix is std_logic_vector(3 downto 0);
	type MemVideoLine is array(0 to DIS_MAX_X - 1) of MemVideoPix;
	type MemVideoFrame is array(0 to DIS_MAX_Y - 1) of MemVideoLine;

	constant VideoFrameA_R : MemVideoFrame:=(
4=>(37|41=>"1100",35|42=>"1101",36=>"1110",others=>"1111"),
5=>(40=>"1101",35=>"1110",others=>"1111"),
6=>(37=>"1101",others=>"1111"),
10=>(34=>"1100",others=>"1111"),
11=>(35=>"1110",others=>"1111"),
12=>(53|54=>"1110",others=>"1111"),
14=>(26=>"1100",48|54=>"1110",others=>"1111"),
15=>(26=>"1100",others=>"1111"),
17=>(41=>"1110",others=>"1111"),
18=>(51=>"1101",40|41|43|48|50=>"1110",others=>"1111"),
19=>(27|39|40|41|43|47=>"1110",others=>"1111"),
20=>(37|38=>"0001",39=>"1010",40=>"1100",41|42|47=>"1110",others=>"1111"),
21=>(36=>"0001",37=>"0010",42=>"0100",41=>"0111",38=>"1001",40|43=>"1101",39|50=>"1110",others=>"1111"),
22=>(36|42|43=>"0100",40|49=>"0101",41=>"1100",37|38|39=>"1110",others=>"1111"),
23=>(47|48=>"0001",49|50=>"0010",39|40|42|43|44=>"0100",41=>"0101",54=>"0111",45=>"1000",30=>"1100",38|55=>"1101",36|37=>"1110",others=>"1111"),
24=>(48|50=>"0001",47|49|54=>"0010",38|53=>"0011",39|41|42|43|44|45|46=>"0100",40=>"0101",25=>"1001",28|31=>"1100",36|37=>"1110",others=>"1111"),
25=>(46|47=>"0000",45|48|49|54|55=>"0001",38|39|40|41|42|43|44|50=>"0100",53=>"1001",25=>"1010",52|56=>"1100",32|33|34|35|36|37=>"1110",others=>"1111"),
26=>(45|46|47|48=>"0000",49|53|54|55=>"0001",39|40|41|42|43|44=>"0100",38|50|51|52|56|57=>"1100",31|32|33|34|35|37=>"1110",others=>"1111"),
27=>(44|45|46|47|55|56|57=>"0000",52|53|54=>"0001",23=>"0010",39|40|41|42|43=>"0100",48=>"0101",49|50|51=>"1100",31|32|33|34|35|36|37|38|58=>"1110",others=>"1111"),
28=>(44|45|46|55|56=>"0000",49|53|54|57=>"0001",47|50|51|52=>"0010",24=>"0011",39|40|41|42|43=>"0100",22=>"0101",58=>"1000",48=>"1100",31|32|33|34|35|36|37|38=>"1110",others=>"1111"),
29=>(44|45|46|47|48|50|51|55|56|57|58=>"0000",49=>"0001",52|53|54=>"0010",38|39|40|41|42|43=>"0100",22=>"1011",30|31|32|33|34|35|36|37|59=>"1110",others=>"1111"),
30=>(44|45|46|47|48|54|55|57|59=>"0000",50|56|58=>"0001",51|52|53=>"0010",27|38|39|40|41|42|43=>"0100",49=>"0101",37=>"0110",25=>"1001",23=>"1101",31|32|33|34|35|36=>"1110",others=>"1111"),
31=>(44|45|46|47|48|55=>"0000",54|56|57|58|59=>"0001",26|49|50|51|52|53=>"0010",37|38|39|40|41|42|43=>"0100",25=>"0110",36=>"1010",27=>"1011",23|24=>"1100",30|31|32|33|34|60=>"1110",others=>"1111"),
32=>(45|46|47=>"0000",44|57|58|59|60=>"0001",25|37|49|50|56=>"0010",26=>"0011",38|39|41|42|43=>"0100",51=>"0101",53|54|55=>"0110",48=>"1000",40|52=>"1001",30|31|32|33|36=>"1110",others=>"1111"),
33=>(44|45|50|51|52|55|56|58|60=>"0000",57|59=>"0001",25|37=>"0010",26=>"0011",36|38|39|41|42|43|53=>"0100",46|54=>"0101",40|49=>"0110",35=>"0111",47|48=>"1010",30=>"1100",21=>"1101",32=>"1110",others=>"1111"),
34=>(50|51|52|54|55|56|57|58|59|60|61=>"0000",53=>"0001",24|25|26|37=>"0010",30|31|38|40|41|42|43=>"0100",39=>"0101",32=>"1000",49=>"1001",44|45|46|47|48=>"1010",27=>"1011",21|35|36=>"1101",20|29|33=>"1110",others=>"1111"),
35=>(50|51|54|55|57|58|59|60|61=>"0000",56=>"0001",24|40|41|43=>"0010",42=>"0100",39=>"0101",20|27|52|53=>"0110",35=>"0111",49=>"1001",44|45|46|47|48=>"1010",29|30|31|37|38=>"1110",others=>"1111"),
36=>(54|55|56|57|58|59|60|61=>"0000",39|43|50=>"0010",40=>"0011",41|42=>"0100",36=>"0111",51|52|53=>"1001",34|44|45|46|47|48|49=>"1010",37|38=>"1100",19|24|27|29=>"1110",others=>"1111"),
37=>(43|54|55|56|57|58|59|60=>"0000",44|50=>"0011",34|41|53|61=>"0100",39|62=>"0101",24|40=>"0110",23|42=>"0111",48|49=>"1000",45|47|51|52=>"1001",46=>"1010",31|35|36|37|38=>"1100",28|29=>"1110",others=>"1111"),
38=>(49|55|56|57|58|60=>"0000",41|52|53|54|59|62=>"0001",38|39=>"0010",35|61=>"0011",50=>"0100",36|51=>"0101",18=>"0111",40=>"1000",47|48=>"1001",44=>"1010",46=>"1011",19|20|23|24|34|37|45=>"1100",28|43=>"1110",others=>"1111"),
39=>(48|49|52|55|56|61=>"0000",38|40|57|60=>"0001",37|53|54|58|59=>"0010",36|51=>"0011",41=>"0100",18|47=>"0101",50=>"1000",46|62=>"1001",19|22|23|26|33|34|35|44|45=>"1100",20=>"1101",27|28|30|42=>"1110",others=>"1111"),
40=>(39|47|48|49|53|54|55|56|58=>"0000",36|37|45|46|51|57|60|61=>"0001",40|52|59=>"0010",62=>"0100",35|38=>"0101",50=>"1001",18|20|21|22|23|33|34=>"1100",19|42=>"1101",27|28|29|41|43|44=>"1110",others=>"1111"),
41=>(35|36|37|38|39|40|43|44|45|46|47|48|49|50|52|53|54|55|57=>"0000",58|60=>"0001",51=>"0010",41=>"0011",32=>"0100",62=>"1000",59=>"1010",34=>"1011",21|33|42|61=>"1100",20=>"1101",22|25|27|28|29|56=>"1110",others=>"1111"),
42=>(37|38|39|41|43|46|49|52|53|54|59|61=>"0000",34|42|45|50|58|60=>"0001",51|55=>"0010",48=>"0100",47=>"0101",44=>"0110",40=>"1000",33=>"1001",57=>"1011",19|20|21|32=>"1100",31|36|62=>"1101",26|27|28|35=>"1110",others=>"1111"),
43=>(42|43|50|51|52|61=>"0000",32|44|59|60=>"0001",40|45|46|49=>"0010",37=>"0011",53|62=>"0110",28=>"0111",47=>"1001",48=>"1011",54=>"1100",17|19|26|27|29|30|31|33|34|35|36|38|39|41=>"1110",others=>"1111"),
44=>(41|42|49|50|51|52=>"0000",62=>"0001",44|45|46=>"0010",48=>"0011",28|31|43|47|53=>"1100",39=>"1101",18|26|27|29|30|32|33|34|35|36|37|38|40=>"1110",others=>"1111"),
45=>(48|49|51|52=>"0000",42|44|50=>"0010",45=>"0100",43|47=>"1000",46=>"1010",27=>"1011",38=>"1100",53=>"1101",28|29|30|31|32|33|34|35|36|37|39|40|54=>"1110",others=>"1111"),
46=>(48|49=>"0000",42=>"0001",47|50|51|52=>"0010",40=>"0101",44|45|46=>"1010",39=>"1100",26|28|29|30|31|32|33|34|35|36|37|38|41=>"1110",others=>"1111"),
47=>(48|49=>"0000",52=>"0001",47|50|51|53|54=>"0010",41=>"0100",43|44|45|46=>"1010",36|37|42=>"1100",29|38|40=>"1101",27|28|30|31|32|33|34|35|39=>"1110",others=>"1111"),
48=>(50|51=>"0000",38|54=>"0001",46|47|48|49|52|53=>"0010",40=>"0011",39=>"0111",45=>"1001",41|42|44|55|56=>"1010",37=>"1011",28|36=>"1100",43=>"1101",24|25|26|27|29|30|31|32|33|34|35=>"1110",others=>"1111"),
49=>(49|50=>"0000",51|52|53|54=>"0001",45|46|47|48=>"0010",55|56=>"0011",44=>"0101",34=>"1000",58=>"1010",37=>"1011",24|38|41=>"1100",25|26|27|28|29|30|32|35|36|39|40=>"1110",others=>"1111"),
50=>(48|50|56=>"0000",43|44|45|49|51|52|53|54|55=>"0001",46|47=>"0010",32=>"1011",36|37|42=>"1100",38=>"1101",25|26|27|29|30|34|35|39|40=>"1110",others=>"1111"),
51=>(48|49|50|55=>"0000",33|43|44|45|51|52|53|54=>"0001",47=>"0010",56=>"0011",37|38=>"1010",36=>"1100",46=>"1101",28|29|31|34|35|39|41|42=>"1110",others=>"1111"),
52=>(47|48|49|50=>"0000",43|45|51|52|53|54=>"0001",44=>"0011",46|56=>"1101",22|26|29|30|32|35|36|55=>"1110",others=>"1111"),
53=>(47|48|49|50=>"0000",51=>"0001",52=>"0111",56=>"1010",46=>"1011",54=>"1101",29|31|33|34|45=>"1110",others=>"1111"),
54=>(57=>"1011",others=>"1111"),
others=>(others=>"1111")
	);
	constant VideoFrameA_G : MemVideoFrame:=(
-- Created Date : 02-Jun-2016 13:29:07
0=>(49=>"1101",others=>"1111"),
1=>(53|54=>"1101",55=>"1110",others=>"1111"),
2=>(52|53=>"1101",others=>"1111"),
3=>(54=>"1100",49|52|53=>"1101",others=>"1111"),
4=>(37|41=>"0001",42=>"0010",35=>"0101",36=>"0111",33=>"1010",38|40=>"1100",39|43=>"1101",44|54=>"1110",others=>"1111"),
5=>(40=>"0010",41=>"0110",35=>"1001",39=>"1010",34|36|37|47|48=>"1011",42=>"1100",33|38|43|44|45|46|49|50|52=>"1101",others=>"1111"),
6=>(37=>"0100",32=>"1001",53=>"1010",33|34|35|36=>"1011",44|45=>"1100",31|38|39|40|41|42|43|46|47|48=>"1101",others=>"1111"),
7=>(50=>"1010",30|32|33|34|35|42=>"1011",43|44|45=>"1100",31|36|37|38|39|40|41|46|47|48|49|52=>"1101",53=>"1110",others=>"1111"),
8=>(31=>"1001",40=>"1010",30|32|33|34|50=>"1011",41|42|43|44|45|46|47|51=>"1100",29|35|36|37|38|39|48|49=>"1101",others=>"1111"),
9=>(28|30=>"0111",29|49=>"1001",48|50=>"1010",31|32|33=>"1011",40|41|42|43|44|45|46|51=>"1100",34|35|36|37|38|39|47=>"1101",52=>"1110",others=>"1111"),
10=>(34=>"0001",32=>"0110",28|45|48=>"1001",49|50|51|54=>"1010",29|30|31|33|35|52=>"1011",38|40|41|42|43|44|46=>"1100",36|37|39|47|53=>"1101",others=>"1111"),
11=>(35=>"0100",27|31|48|51=>"1001",36|50=>"1010",29|30|32|33|34|47|53=>"1011",41|42|43|44|45|46=>"1100",28|37|38|39|40|49|52=>"1101",others=>"1111"),
12=>(53=>"0100",35=>"0101",30|34=>"0110",51=>"0111",29|36|43|54=>"1000",25|27|33=>"1001",31|46|47|50|52=>"1010",26|28|32|44=>"1011",40|41|42|45|48=>"1100",37|38|39|49=>"1101",others=>"1111"),
13=>(34|35|37=>"0101",33=>"0110",28|36=>"0111",45|54=>"1000",30|31|32|46|47|52|53=>"1001",50|51=>"1010",29|40|43=>"1011",27|38|39|41|42|44|48=>"1100",26|49=>"1101",others=>"1111"),
14=>(26=>"0001",54=>"0100",34|35|37=>"0101",29|32|33=>"0110",41=>"1000",30|31|38|51=>"1001",27|48|49|50|53=>"1010",28=>"1011",36|39|40|42|43|44|45|46|47=>"1100",25|52=>"1101",others=>"1111"),
15=>(26=>"0010",29|34|36=>"0101",28|30|31|32|33|37|38=>"0110",27|35|41=>"1000",42|44|50|53=>"1001",48|49|51|55=>"1010",43=>"1011",39|40|45|46|47|52|54=>"1100",25=>"1101",others=>"1111"),
16=>(30|31|33|35|36|38=>"0101",32=>"0110",29=>"0111",28|34|41=>"1000",46|48|49|50=>"1001",25|37|42|43|44|45|47|51|52|53|54|55=>"1010",26|40=>"1011",39=>"1100",27=>"1101",others=>"1111"),
17=>(41=>"0001",30|31|32|33|34|35|39=>"0101",37=>"0110",29=>"0111",27|44|45|46|47|48=>"1000",25|28|42=>"1001",26|43|52|54|55=>"1010",36|40|53=>"1011",38|49|50|51=>"1100",24=>"1101",others=>"1111"),
18=>(41|48=>"0001",40=>"0010",43=>"0011",32|33|36|37|38=>"0101",24|29=>"0110",28|30|31|35=>"0111",26|42|47=>"1000",27|45=>"1001",25|34|44|46|49|51|52|53=>"1010",54=>"1011",39|50|55=>"1100",56=>"1110",others=>"1111"),
19=>(39|40|41|47=>"0001",43=>"0100",33|34|35|37=>"0101",27|28|29|30|31|32=>"0111",36=>"1000",25|26|38|48=>"1001",46|49|50|51|52|53|54|55=>"1010",42|44|45=>"1100",24=>"1101",others=>"1111"),
20=>(40|41|42=>"0001",37|38|47=>"0010",34|35=>"0101",33=>"0110",24|28|29|30|31|32|39=>"0111",27|36|44|51|52=>"1000",26|48=>"1001",25|49|50|53|54|55=>"1010",56=>"1011",43|45|46=>"1100",others=>"1111"),
21=>(38|39|40|43=>"0001",36|37|41=>"0010",42=>"0011",33|34=>"0101",35=>"0110",24|28|29|30|31|32=>"0111",26|27|44|45|46|47|51=>"1000",25|48|49|52=>"1001",50|53|54|55=>"1010",56=>"1101",others=>"1111"),
22=>(37|38|39=>"0001",36|40=>"0011",42|43|49=>"0100",33|35=>"0101",26|27|28|30|31|32|34|41=>"0111",24|51=>"1000",29|48=>"1001",44|45|46|47|55|56=>"1010",50|52|54=>"1100",25|53=>"1101",others=>"1111"),
23=>(30|36|37|38=>"0001",48=>"0010",49|50=>"0011",39|40|41|42|43|44=>"0100",32|33|34|35|45=>"0101",26|27|29|31=>"0111",28|51|54=>"1001",46|52|55|56=>"1010",25|53=>"1100",24=>"1101",47=>"1110",others=>"1111"),
24=>(28|31|36|37=>"0001",38|50=>"0010",49=>"0011",35|39|40|41|42|43|44|45=>"0100",25|32|33|34|46=>"0101",27=>"0110",26|29|30=>"0111",53|54=>"1000",47|48=>"1001",55|56=>"1010",24|51|52=>"1101",others=>"1111"),
25=>(32|33|34|35|36|37|52|53|56=>"0001",55=>"0010",38=>"0011",25|39|40|41|42|43|44|50=>"0100",26|31=>"0110",27|29|30|54=>"0111",28|49=>"1000",45|46|47=>"1010",24|51=>"1101",23|48=>"1110",others=>"1111"),
26=>(31|32|37|50|51|52|56=>"0001",33|34|35|36|38|49|54|55=>"0010",39|40|41|42|43|44=>"0100",25|26|27=>"0110",28|29|30|53=>"0111",23|45|47=>"1010",24=>"1101",46|48|57=>"1110",others=>"1111"),
27=>(50|51=>"0001",31|32|33|34|35|36|37|38|54=>"0010",23=>"0011",39|40|41|42|43=>"0100",24|25|26|55=>"0110",27|28|29|30|52|53=>"0111",56|57=>"1000",44|45|47=>"1010",48=>"1100",22=>"1101",46|49=>"1110",others=>"1111"),
28=>(38=>"0001",24|31|32|33|34|35|36|37|49|54=>"0010",47|57=>"0011",22|39|40|41|42|43|53=>"0100",26=>"0110",27|28|29|30|52=>"0111",50|51|55|56=>"1000",25|58=>"1001",23|44|45|46=>"1010",48=>"1110",others=>"1111"),
29=>(30|31|32|33|34|35|36|37=>"0010",58=>"0011",38|39|40|41|42|43|49=>"0100",24|25|54|57=>"0110",22|23|26|27|28|29|53=>"0111",55|56=>"1000",44|45|46|48|52=>"1010",47=>"1011",50|51=>"1101",others=>"1111"),
30=>(31|32|33|34|35|36|56=>"0010",27|37|38|39|40|41|42|43|58=>"0100",23|25=>"0101",29|49|54=>"0110",26|28|30=>"0111",51|52|53|55|57=>"1000",22|44|45|47|48|59=>"1010",50=>"1100",21|24|46=>"1101",others=>"1111"),
31=>(23|24=>"0001",25|30|31|32|33|34|36|54|58=>"0010",26|37|38|39|40|41|42|43=>"0100",28|59=>"0101",29|35|56|57=>"0110",27|49|50|52|53=>"1000",51=>"1001",44|45|46|47|48=>"1010",21|22=>"1101",20|55=>"1110",others=>"1111"),
32=>(30|31|32|33|60=>"0010",25|37=>"0011",26|38|39|40|41|42|43=>"0100",58|59=>"0101",57=>"0110",24|28|29|34|35|50=>"0111",49|56=>"1000",44|48=>"1001",20|23|27|36|45|46|47|51|55=>"1010",52|53|54=>"1011",21=>"1100",22=>"1101",others=>"1111"),
33=>(21=>"0001",30|32|53=>"0010",25|26|37=>"0011",36|38|39|40|41|42|43=>"0100",27|35|58|59|60=>"0101",33|57=>"0110",22|23|24=>"0111",28|54=>"1000",49|50|52=>"1001",34|44|45|51|55=>"1010",29|31|46=>"1011",20|47|48=>"1100",19|56=>"1110",others=>"1111"),
34=>(35|36=>"0001",53=>"0010",21|24|25|26|37=>"0011",30|31|33|38|39|40|41|42|43|60=>"0100",20|27|32|57=>"0101",28|56=>"0110",22|23|34|58=>"0111",19|54|55|59|61=>"1000",29|50|51=>"1010",44|45|46|47|48|49|52=>"1100",others=>"1111"),
35=>(37|38=>"0001",27|30=>"0010",20|24|29|40|41|43=>"0011",35|39|42|59=>"0100",60=>"0101",34|36=>"0110",19|22|23|28|31|32|33=>"0111",51|54|57|58|61=>"1000",21=>"1001",25|26|50|52=>"1010",53=>"1011",44|45|46|47|48|49=>"1100",18|55|56=>"1110",others=>"1111"),
36=>(37|38=>"0001",27|28|29=>"0010",26|36=>"0011",39|40|41|42=>"0100",20|21|22|23|59=>"0101",34|35=>"0110",30|31|32|33=>"0111",56|57|58|60|61=>"1000",19|24|50|54=>"1001",25|43=>"1010",51|52|53=>"1011",44|45|46|47|48|49=>"1100",18=>"1101",55=>"1110",others=>"1111"),
37=>(31|35|36|37|38=>"0001",28|29|61=>"0010",39|44=>"0011",20|23|34|40|41|42=>"0100",19|21|22|24|25|27=>"0101",30=>"0110",26|32|33=>"0111",57|58|59|60=>"1000",53|55|56=>"1001",43=>"1010",47|48|49|51|52|62=>"1011",18|45|46=>"1100",50=>"1101",54=>"1110",others=>"1111"),
38=>(18|19|20|23|24|34|37=>"0001",27|28|36|41=>"0010",61=>"0011",26|35|38|39|40|44|58=>"0100",21|25|59=>"0101",29|42|43|53|54=>"0110",30|31|32|33=>"0111",49=>"1000",55|56|57=>"1001",60=>"1010",47|48=>"1011",22|50|51|62=>"1100",46=>"1101",45|52=>"1110",others=>"1111"),
39=>(19|22|23|26|33|34|35|62=>"0001",27|28|30|38|40|41=>"0010",18|20|36=>"0011",37=>"0100",24|29|42|43|60=>"0101",39|53|54|57|58|59=>"0110",25|31|32|47=>"0111",56=>"1000",48=>"1001",21=>"1010",46|49|50=>"1011",51=>"1101",44|45|52|55|61=>"1110",others=>"1111"),
40=>(18|20|21|22|23|33|34|35=>"0001",19|25|26|27|29|36|37|45|46=>"0010",38=>"0011",42=>"0100",28|41|43|44|60|61=>"0101",24|52|59|62=>"0110",30|31|32|40|55|56=>"0111",39|47|48|49|58=>"1001",57=>"1010",50=>"1011",51|53=>"1101",54=>"1110",others=>"1111"),
41=>(21|33|34|59=>"0001",25|27|28|29|32|61=>"0010",20=>"0011",35|60=>"0101",31|51=>"0110",22|30=>"0111",58=>"1000",18|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|54|55|57=>"1001",62=>"1011",19|23|26=>"1100",52|53=>"1110",others=>"1111"),
42=>(19|20|21|32|33=>"0001",26|27|28|31|34|35|36=>"0010",54=>"0100",60=>"0101",22|30|50|51|58=>"0110",29|40|45=>"0111",48=>"1000",37|38|39|41|42|43|46|49|59=>"1001",61=>"1010",44|47|55=>"1011",18=>"1100",25|53|57=>"1101",52|62=>"1110",others=>"1111"),
43=>(33|34|35|36=>"0001",26|27|32|37=>"0010",28=>"0011",29|30|31|51=>"0100",38|39|41|50|59|60=>"0101",46|49=>"0110",40|44|45=>"0111",42|43|53|62=>"1001",61=>"1010",17|19=>"1011",20|47=>"1100",25=>"1101",21|48|52|54=>"1110",others=>"1111"),
44=>(31|32|33|34|35|36=>"0001",26|28=>"0010",39=>"0011",27|29|30|49|51=>"0100",37|38|40|62=>"0101",44=>"0110",45|46|48|50=>"0111",18|43=>"1000",41|42|52=>"1001",47|53=>"1110",others=>"1111"),
45=>(27|32|33|34|35|38=>"0001",30|31|36=>"0010",29=>"0100",37|39|40|41=>"0101",28=>"0110",42|44=>"0111",50=>"1000",43|45=>"1001",47|48|49|51|52=>"1010",46=>"1100",others=>"1111"),
46=>(32|33|34|39=>"0001",29|30|31|35|40=>"0010",28|38=>"0100",26|36|37=>"0101",41|42=>"0110",47|50|52=>"1000",51=>"1001",48|49=>"1010",43=>"1011",44|45|46=>"1100",others=>"1111"),
47=>(29|31|32|33|34|36|37|41=>"0001",30|38|40=>"0010",27|28|39=>"0100",35=>"0101",26|47|50|51|53|54=>"1000",48|49|52=>"1010",42|43|44|45|46=>"1100",25=>"1101",others=>"1111"),
48=>(28|30|31|32|33|34|35|36|39=>"0001",37|38|40=>"0010",25|26|27=>"0100",24=>"0101",54=>"0110",46|47|49|52|53=>"1000",29|48=>"1001",50|51=>"1010",45|55=>"1011",41|42|43|44|56=>"1100",others=>"1111"),
49=>(29|30|35|36|37|38|39=>"0001",24|32|54=>"0010",25|26|27|56=>"0100",28|31=>"0101",40|43|52|53=>"0110",34|45=>"0111",44|46|47|48|55=>"1000",33|41|49|50|51|58=>"1010",42=>"1011",23=>"1101",others=>"1111"),
50=>(29|30|34|35|36|37|38|39=>"0001",40|43|44|53|54=>"0010",26|27=>"0100",25|41|51|52|55|56=>"0110",28|45|46|47=>"0111",49=>"1001",31|33|42|48|50=>"1010",24|32=>"1100",22|23=>"1110",others=>"1111"),
51=>(29|30|31|34|35|36|38=>"0001",28|37|39|43|44|52|53=>"0010",25=>"0101",40|41|42|45|51|54=>"0110",47|49|55=>"0111",26|27=>"1001",46|48|50=>"1010",23|24|32|56=>"1100",33=>"1101",others=>"1111"),
52=>(36=>"0001",30|32|43|51|52=>"0010",29=>"0100",22|26|34|35=>"0101",28|44|45|53|54=>"0110",49=>"1000",25|27|47|48|50=>"1010",46=>"1011",24|31|33|37=>"1100",55=>"1110",others=>"1111"),
53=>(33=>"0001",29|31|34|51=>"0010",32=>"0111",49|50=>"1000",28|52=>"1001",47|48=>"1010",30=>"1100",35|45|46|56=>"1110",others=>"1111"),
54=>(57=>"1101",others=>"1111"),
55=>(27|28=>"1010",23|24=>"1110",others=>"1111"),
56=>(26=>"1010",24=>"1100",20=>"1101",others=>"1111"),
57=>(23=>"0100",others=>"1111"),
others=>(others=>"1111")
	);
	constant VideoFrameA_B : MemVideoFrame:=(
-- Created Date : 02-Jun-2016 13:29:38
0=>(49=>"0101",others=>"1111"),
1=>(53=>"0100",54=>"0101",55=>"1100",51=>"1110",others=>"1111"),
2=>(52|53=>"0100",49=>"1100",others=>"1111"),
3=>(49|52|53=>"0100",48=>"1110",others=>"1111"),
4=>(40=>"0110",43=>"1000",44=>"1010",56=>"1011",33|38=>"1100",36|39|45|52=>"1101",42=>"1110",others=>"1111"),
5=>(47=>"0011",48|49|50|52=>"0100",44|45=>"0101",43=>"0110",41=>"0111",46=>"1011",34|36|37|42=>"1100",33|35|38|39|40=>"1101",others=>"1111"),
6=>(45|46|47|48=>"0100",44=>"0101",41|42|43=>"0110",39=>"1000",40=>"1011",32|33|34|35|36=>"1100",38=>"1101",31|53=>"1110",others=>"1111"),
7=>(50=>"0010",45|48=>"0011",42|46|47|52=>"0100",43|44=>"0101",40|41=>"0110",49=>"1000",33|34|35|39=>"1100",31|32|36|37|38=>"1101",30=>"1110",others=>"1111"),
8=>(40|50=>"0010",46|47|48|49|51=>"0011",44|45=>"0100",41|42|43=>"0101",39=>"0110",31=>"1001",37=>"1010",38|52=>"1011",32|33|34=>"1100",29|30|35|36=>"1101",others=>"1111"),
9=>(49|50=>"0001",48=>"0010",46|47|51=>"0011",43|44|45=>"0100",40|41|42=>"0101",30=>"0110",52=>"1010",28=>"1011",29|31|32|33|38|39=>"1100",34|35|36|37=>"1101",others=>"1111"),
10=>(48=>"0001",45|50|51|52=>"0010",46|47|49|54=>"0011",32|41|42|43|44=>"0100",40=>"0101",38=>"0111",37=>"1000",53=>"1010",28|29|30|31|33|35=>"1100",36|39=>"1101",others=>"1111"),
11=>(48|51=>"0001",47|50=>"0010",46|49|52=>"0011",42|43|44|45|53=>"0100",41=>"0101",31|36=>"1001",35=>"1010",27|29|30|32|33|34|39=>"1100",28|37|38|40=>"1101",others=>"1111"),
12=>(36|43|50|52=>"0010",44|47|48|49=>"0011",35|40|41|42|45|46=>"0100",30|34|51=>"0101",29=>"0111",53|54=>"1011",25|27|28|31|32|33=>"1100",26|37|38|39=>"1101",others=>"1111"),
13=>(52|53=>"0001",45|47|50|51=>"0010",40|42|43|48|49=>"0011",34|35|36|39|41|44|46|54=>"0100",28=>"0101",37=>"1001",31|33=>"1011",27|29|30|32|38=>"1100",26=>"1101",others=>"1111"),
14=>(51=>"0001",41|49|50|53=>"0010",42|47|48|52=>"0011",34|35|36|39|40|43|44|45|46=>"0100",29=>"0101",37=>"0111",38=>"1001",32|33|54=>"1011",27|28|30|31=>"1100",25=>"1101",55=>"1110",others=>"1111"),
15=>(50|53=>"0001",41|43|44|48|49|51|55=>"0010",35|52|54=>"0011",29|34|36|37|38|39|40|42|45|46|47=>"0100",30=>"0101",27=>"0111",33=>"1010",28|31|32=>"1011",25=>"1101",others=>"1111"),
16=>(49|50=>"0001",34|41|51|52|53|54|55=>"0010",37=>"0011",30|33|35|36|38|39|40|42|43|44|45|46|47|48=>"0100",31=>"0101",29=>"0110",32=>"1011",25|26|28=>"1100",27=>"1101",others=>"1111"),
17=>(44|45|46|47|48|54|55=>"0010",42|49|53=>"0011",30|31|33|34|35|36|37|38|40|43|50|51|52=>"0100",29|32=>"0110",39=>"0111",27|28=>"1011",25|26=>"1100",24=>"1101",41=>"1110",others=>"1111"),
18=>(42|45|47=>"0010",35|44|46|49|54|55=>"0011",32|33|34|36|37|39|50|52|53=>"0100",29|30|31|38|51=>"0101",28=>"0110",26=>"0111",24|56=>"1011",25|27|43=>"1100",40|48=>"1110",others=>"1111"),
19=>(48|53|54|55=>"0010",36|37|49=>"0011",33|34|35|42|44|45|50|51|52=>"0100",28|29|30|31|32|38|46=>"0101",27|43=>"1010",25|26=>"1100",24=>"1101",40|56=>"1110",others=>"1111"),
20=>(44|51|52|54=>"0010",33|34|35|48|53|55|56=>"0011",36|43|45|46|49|50=>"0100",28|29|30|31|32|39=>"0101",37|38=>"0110",24=>"0111",25|26|27=>"1100",40|47=>"1101",others=>"1111"),
21=>(44|45|46|47|51|52|53|54=>"0010",34|35|55=>"0011",33|48|49|50=>"0100",28|29|30|31|32=>"0101",24|36|37=>"0110",56=>"1000",42=>"1001",27=>"1010",26|41=>"1011",25|38=>"1100",others=>"1111"),
22=>(34|44|45|48|51|55|56=>"0010",33|35|46|47=>"0011",50|54=>"0100",28|30|31|32|52=>"0101",36|53=>"0110",24|27|49=>"0111",40=>"1001",29|42|43=>"1010",26|41=>"1011",25=>"1101",others=>"1111"),
23=>(46|51|52|56=>"0010",33|34|35=>"0011",32|55=>"0100",29|31|53=>"0101",26|27|48=>"0110",37|50=>"0111",39|40=>"1000",45|49|54=>"1001",28|41|42|43|44=>"1010",24|25=>"1101",others=>"1111"),
24=>(55|56=>"0010",33|34=>"0011",32|35=>"0100",29|30=>"0101",26|51|52=>"0110",36|37|38|50=>"0111",39=>"1000",25|27|49=>"1001",40|41|42|43|44|45|46=>"1010",47|48|53|54=>"1100",24=>"1101",others=>"1111"),
25=>(31=>"0100",29|30|51|55=>"0110",28|32|33|34|35|36|37=>"0111",38=>"1000",25|50=>"1001",27|39|40|41|42|43|44=>"1010",26|49=>"1011",45|53|54=>"1100",24|46|47=>"1101",23=>"1110",others=>"1111"),
26=>(28|29|30|49|54=>"0110",31|32|37|38|55=>"0111",36=>"1000",33|34|35=>"1001",23|39|40|41|42|43|44=>"1010",25|26|27=>"1011",53=>"1100",24|45|47=>"1101",57=>"1110",others=>"1111"),
27=>(27|28|29|30|54=>"0110",23=>"0111",31=>"1000",32|33|34|35|36|37|38=>"1001",39|40|41|42|43|55=>"1010",24|25|26=>"1011",52|53|56|57=>"1100",44|45|47|48=>"1101",49=>"1110",others=>"1111"),
28=>(27|28|29|30|54=>"0110",24|49=>"0111",22|57=>"1000",31|32|33|34|35|36|37|47|53=>"1001",23|25|39|40|41|42|43=>"1010",26=>"1011",50|51|52|55|56|58=>"1100",44|45|46=>"1101",48=>"1110",others=>"1111"),
29=>(23|26|27|28|29=>"0110",58=>"0111",49=>"1000",30|31|32|33|34|35|36|37=>"1001",24|38|39|40|41|42|43|57=>"1010",22|25=>"1011",48|53|54|55|56=>"1100",44|45|46|47|52=>"1101",others=>"1111"),
30=>(26|29|30|56=>"0110",25|28=>"0111",27|58=>"1000",31|32|33|34|35|36=>"1001",22|37|38|39|40|41|42|43|49|54=>"1010",51|52|53|55|57|59=>"1100",21|24|44|45|47|48=>"1101",46|50=>"1110",others=>"1111"),
31=>(28=>"0100",29=>"0110",54|58=>"0111",26|30|31|32|33|34|36=>"1001",27|35|37|38|39|40|41|42|43|59=>"1010",56|57=>"1011",25|49|50|51|52|53=>"1100",20|21|22|44|45|46|47|48=>"1101",others=>"1111"),
32=>(34|35=>"0101",28|29=>"0110",24|60=>"0111",30=>"1000",25|26|31|32|33|37=>"1001",23|27|38|39|40|41|42|43|58|59=>"1010",20|48|50|57=>"1011",21|36|44|49|51|53|54|55|56=>"1100",22|45|46|47|52=>"1101",others=>"1111"),
33=>(27=>"0100",22|23|24|33=>"0110",28=>"0111",53=>"1000",25|26|30|32|35|37|60=>"1001",34|36|38|39|40|41|42|43|58|59=>"1010",49|54|57=>"1011",20|29|31|44|46|50|52|55=>"1100",19|45|47|48|51=>"1101",others=>"1111"),
34=>(34=>"0101",22|23|27|28=>"0110",19|53=>"0111",20|24|25|26|32|37|60=>"1001",30|31|38|40|41|42|43|56|57=>"1010",39|58=>"1011",29|33|54|55|59|61=>"1100",44|45|46|47|48|49|50|51=>"1101",21|52=>"1110",others=>"1111"),
35=>(33=>"0101",22|23|28|31|32=>"0110",19|20=>"0111",27=>"1000",24|29|30|34|40|41|43|59=>"1001",21|25|26|39|42|60=>"1010",35|36=>"1011",51|52|53|54|57|58|61=>"1100",44|45|46|47|48|49|50=>"1101",18=>"1110",others=>"1111"),
36=>(20|21|22|23=>"0100",26|30|31|32|33=>"0110",18=>"0111",34=>"1000",27|28|29|39|40=>"1001",24|25|41|42|59=>"1010",35|50=>"1011",19|36|43|51|52|53|54|56|57|58|60|61=>"1100",44|45|46|47|48|49=>"1101",others=>"1111"),
37=>(19|21|22|25=>"0100",18=>"0101",20|26|32|33=>"0110",23|27|30|44=>"0111",42=>"1000",24|28|29=>"1001",34|39|41=>"1010",40|55|56|60|61=>"1011",47|48|49|51|52|53|57|58|59=>"1100",43|45|46|62=>"1101",50=>"1110",others=>"1111"),
38=>(21|25=>"0100",22=>"0101",29|30|31|32|33|41=>"0110",26=>"0111",44=>"1000",27|28|35|38|39|58=>"1001",40|43|53|54|59=>"1010",18|36|42|49|55|56|57|61=>"1011",47|48|60=>"1100",46|51|62=>"1101",45|50=>"1110",others=>"1111"),
39=>(24=>"0100",18|25|31|32|40=>"0110",21|29|41=>"0111",38=>"1000",27|28|30|36|37|42|43|60=>"1001",47|53|54|57|58|59=>"1010",39|48|56=>"1011",20|46|50=>"1100",49=>"1101",44|45|51|62=>"1110",others=>"1111"),
40=>(24=>"0101",30|31|32|36|37|45|46=>"0110",38=>"0111",25=>"1000",26|27|29|41|42|43|44=>"1001",28|35|40|52|59|60|61=>"1010",39|47|48|49|55|56|58|62=>"1011",50|57=>"1100",19|53=>"1110",others=>"1111"),
41=>(18=>"0011",19|23=>"0101",26|30=>"0110",25|27|28|29|35=>"1001",22|32|51|60=>"1010",31|36|37|38|39|40|41|43|44|45|46|47|48|49|50|54|57|58=>"1011",42|55|62=>"1100",20=>"1101",34|59=>"1110",others=>"1111"),
42=>(22=>"0100",18=>"0101",25|29=>"0110",34|35|36=>"0111",26|27|28|54=>"1001",50|51|58|60=>"1010",30|37|38|39|40|41|42|43|45|46|48|49=>"1011",44|47|59|61=>"1100",33|55=>"1101",31|57|62=>"1110",others=>"1111"),
43=>(20=>"0101",19|32=>"0110",33|35|36|37=>"0111",28=>"1000",26|27|34|41|50|51=>"1001",29|39|46|49|59|60=>"1010",30|31|42|44|45|53=>"1011",21|38|40|43|61|62=>"1100",47=>"1101",25|48|54=>"1110",others=>"1111"),
44=>(32|33|34|35|36=>"0111",26|49|51=>"1001",29|44|62=>"1010",27|30|41|42|43|45|46|48|50|52=>"1011",37|38|40=>"1100",53=>"1101",18|28|39|47=>"1110",others=>"1111"),
45=>(32|33|34|35=>"0111",36=>"1000",30|31|41=>"1001",28|29|42|44=>"1011",37|39|40|43|45|47|50=>"1100",46|48|49|51|52=>"1101",53=>"1110",others=>"1111"),
46=>(32|33|34|35=>"0111",29|30|31|36|38=>"1001",28|37=>"1010",26|40|41|42=>"1011",47|50|51|52=>"1100",44|45|46|48|49=>"1101",43=>"1110",others=>"1111"),
47=>(31|32|33|34=>"0111",30|35|41=>"1001",28|29|39=>"1010",27=>"1011",26|47|49|50|51|52|53|54=>"1100",38|42|43|44|45|46|48=>"1101",25|40=>"1110",others=>"1111"),
48=>(38=>"0110",30|31|32|33|34|37=>"0111",35|40=>"1000",26=>"1010",24|25|27|29|54=>"1011",39|45|46|47|48|49|52|53=>"1100",41|42|43|44|50|51|55=>"1101",56=>"1110",others=>"1111"),
49=>(33=>"0101",29|30|32|35|36|39|54=>"0111",28|31|56=>"1001",25=>"1010",26|27|34|40|43|44|45|52|53|55=>"1011",41|46|47|48|51|58=>"1100",24|49|50=>"1101",42=>"1110",others=>"1111"),
50=>(24|33=>"0101",44|53=>"0110",29|30|34|35|39|43|54=>"0111",32=>"1000",25|40=>"1001",27|28|31|55|56=>"1010",26|41|45|46|47|51|52=>"1011",38|42|48|49=>"1100",23|50=>"1101",22=>"1110",others=>"1111"),
51=>(23|24|32=>"0101",43|44=>"0110",28|29|30|31|34|35|37|52|53=>"0111",25|39=>"1001",26|27=>"1010",40|41|42|45|47|49|51|54|55=>"1011",50=>"1100",46|48=>"1101",38|56=>"1110",others=>"1111"),
52=>(31|33=>"0101",51|52=>"0110",30|32|36|43=>"0111",26|28|29|35=>"1001",27|34|44=>"1010",22|45|53|54=>"1011",25|49|50=>"1100",24|37|46|47|48=>"1101",others=>"1111"),
53=>(30=>"0101",28|32=>"0110",29|31|33|34|51=>"0111",49|50|52=>"1011",47|48=>"1101",35|56=>"1110",others=>"1111"),
54=>(57=>"1101",22=>"1110",others=>"1111"),
55=>(27=>"1010",28=>"1011",23=>"1101",24=>"1110",others=>"1111"),
56=>(26=>"1010",20|24=>"1101",others=>"1111"),
57=>(23=>"1001",others=>"1111"),
others=>(others=>"1111")
	);
end package;