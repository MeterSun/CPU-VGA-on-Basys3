-- Created Date : 06-Jun-2016 12:10:23
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use work.comMCU.AlL;
package HEXfile is
	constant ROM:MEMORY:=(
X"75",X"C7",X"00",X"75",X"C8",X"58",X"75",X"C9",X"23",X"75",X"C6",X"FF",X"75",X"A0",X"F5",X"75",
X"B0",X"0F",X"75",X"20",X"FF",X"75",X"20",X"00",X"75",X"A0",X"F6",X"75",X"B0",X"0F",X"75",X"20",
X"FF",X"75",X"20",X"00",X"75",X"A0",X"F7",X"75",X"B0",X"08",X"75",X"20",X"FF",X"75",X"20",X"00",
X"75",X"80",X"00",X"75",X"80",X"11",X"75",X"A0",X"F0",X"75",X"B0",X"00",X"75",X"20",X"FF",X"75",
X"20",X"00",X"7F",X"08",X"7E",X"FF",X"7D",X"FF",X"DD",X"FE",X"DE",X"FA",X"DF",X"F6",X"75",X"80",
X"10",X"75",X"A0",X"F0",X"75",X"B0",X"01",X"75",X"20",X"FF",X"75",X"20",X"00",X"7F",X"08",X"7E",
X"FF",X"7D",X"FF",X"DD",X"FE",X"DE",X"FA",X"DF",X"F6",X"75",X"A0",X"F0",X"75",X"B0",X"02",X"75",
X"20",X"FF",X"75",X"20",X"00",X"75",X"A0",X"E0",X"75",X"B0",X"30",X"75",X"20",X"FF",X"75",X"20",
X"00",X"75",X"A0",X"E1",X"75",X"B0",X"31",X"75",X"20",X"FF",X"75",X"20",X"00",X"75",X"A0",X"E2",
X"75",X"B0",X"32",X"75",X"20",X"FF",X"75",X"20",X"00",X"75",X"A0",X"E3",X"75",X"B0",X"33",X"75",
X"20",X"FF",X"75",X"20",X"00",X"75",X"A0",X"E4",X"75",X"B0",X"34",X"75",X"20",X"FF",X"75",X"20",
X"00",X"75",X"A0",X"E5",X"75",X"B0",X"35",X"75",X"20",X"FF",X"75",X"20",X"00",X"75",X"A0",X"E6",
X"75",X"B0",X"36",X"75",X"20",X"FF",X"75",X"20",X"00",X"75",X"A0",X"E7",X"75",X"B0",X"37",X"75",
X"20",X"FF",X"75",X"20",X"00",X"75",X"A0",X"E8",X"75",X"B0",X"38",X"75",X"20",X"FF",X"75",X"20",
X"00",X"75",X"A0",X"E9",X"75",X"B0",X"39",X"75",X"20",X"FF",X"75",X"20",X"00",X"7F",X"0F",X"7E",
X"FF",X"7D",X"FF",X"DD",X"FE",X"DE",X"FA",X"DF",X"F6",X"75",X"A0",X"E0",X"85",X"CF",X"B0",X"75",
X"20",X"FF",X"75",X"20",X"00",X"75",X"A0",X"E1",X"85",X"CE",X"B0",X"75",X"20",X"FF",X"75",X"20",
X"00",X"75",X"A0",X"E2",X"85",X"CD",X"B0",X"75",X"20",X"FF",X"75",X"20",X"00",X"75",X"A0",X"E3",
X"85",X"CC",X"B0",X"75",X"20",X"FF",X"75",X"20",X"00",X"75",X"A0",X"E8",X"85",X"CB",X"B0",X"75",
X"20",X"FF",X"75",X"20",X"00",X"75",X"A0",X"E9",X"85",X"CA",X"B0",X"75",X"20",X"FF",X"75",X"20",
X"00",X"75",X"A0",X"E4",X"85",X"C1",X"B0",X"75",X"20",X"FF",X"75",X"20",X"00",X"75",X"A0",X"E5",
X"75",X"B0",X"00",X"75",X"20",X"FF",X"75",X"20",X"00",X"75",X"A0",X"E6",X"75",X"B0",X"00",X"75",
X"20",X"FF",X"75",X"20",X"00",X"75",X"A0",X"E7",X"75",X"B0",X"00",X"75",X"20",X"FF",X"75",X"20",
X"00",X"85",X"C1",X"90",X"A8",X"C0",X"B8",X"5A",X"17",X"85",X"C3",X"A0",X"85",X"C2",X"B0",X"75",
X"20",X"FF",X"75",X"20",X"00",X"75",X"90",X"FF",X"7E",X"FF",X"7D",X"FF",X"DD",X"FE",X"DE",X"FA",
X"02",X"00",X"F9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
X"00");
end;
